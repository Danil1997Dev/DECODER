// SysFiltr_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module SysFiltr_tb #(parameter
CLK_PRD = 20,
T_100=50_000_000/50_000_000, 
N_100=50_000_000/440_000,
T_50=50_000_000/25_000_000, 
N_50=25_000_000/440_000,
T_5=50_000_000/5_000_000, 
N_5=5_000_000/440_000,
K=350)(); 
	logic [31:0] signal_100_i,signal_50_i,signal_5_i;
	logic indicate_100,indicate_50,indicate_5;
	logic work_100 = 1;
	logic work_50 = 1;
	logic work_5 = 1;

	logic [31:0] mem_100_a [0:K*N_100-1];  
	logic [31:0] mem_100_b [0:K*N_100-1];
	logic [31:0] mem_100_c [0:K*N_100-1]; 

	logic [31:0] mem_50_a [0:K*N_50-1];  
	logic [31:0] mem_50_b [0:K*N_50-1];
	logic [31:0] mem_50_c [0:K*N_50-1]; 

	logic [31:0] mem_5_a [0:K*N_5-1];  
	logic [31:0] mem_5_b [0:K*N_5-1];
	logic [31:0] mem_5_c [0:K*N_5-1]; 

	logic sysfiltr_inst_clk_bfm_clk_clk;       // SysFiltr_inst_clk_bfm:clk -> [SysFiltr_inst:clk_clk, SysFiltr_inst_reset_bfm:clk]
	logic sysfiltr_inst_reset_bfm_reset_reset; // SysFiltr_inst_reset_bfm:reset -> SysFiltr_inst:reset_reset_n

	SysFiltr #(.CLK_REF(50_000_000),.SAMPL_T(50_000_000),.FRQ_SIGNAL(440_000),.FRQ_DELT(44_000)) sysfiltr_100_inst (
		.clk_clk                 (sysfiltr_inst_clk_bfm_clk_clk),       //            clk.clk 
		.decoder_expend_signal_i (signal_100_i),                                    //               .signal_i
		.decoder_expend_work (work_100),                                    //               .work
		.decoder_expend_indicate (indicate_100),                                    //               .indicate
		.reset_reset_n           (sysfiltr_inst_reset_bfm_reset_reset)  //          reset.reset_n
	);

	SysFiltr #(.CLK_REF(50_000_000),.SAMPL_T(25_000_000),.FRQ_SIGNAL(440_000),.FRQ_DELT(44_000)) sysfiltr_50_inst (
		.clk_clk                 (sysfiltr_inst_clk_bfm_clk_clk),       //            clk.clk 
		.decoder_expend_signal_i (signal_50_i),                                    //               .signal_i
		.decoder_expend_work (work_50),                                    //               .work
		.decoder_expend_indicate (indicate_50),                                    //               .indicate
		.reset_reset_n           (sysfiltr_inst_reset_bfm_reset_reset)  //          reset.reset_n
	);

	SysFiltr #(.CLK_REF(50_000_000),.SAMPL_T(5_000_000),.FRQ_SIGNAL(440_000),.FRQ_DELT(44_000)) sysfiltr_5_inst (
		.clk_clk                 (sysfiltr_inst_clk_bfm_clk_clk),       //            clk.clk 
		.decoder_expend_signal_i (signal_5_i),                                    //               .signal_i
		.decoder_expend_work (work_5),                                    //               .work
		.decoder_expend_indicate (indicate_5),                                    //               .indicate
		.reset_reset_n           (sysfiltr_inst_reset_bfm_reset_reset)  //          reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sysfiltr_inst_clk_bfm (
		.clk (sysfiltr_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) sysfiltr_inst_reset_bfm (
		.reset (sysfiltr_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (sysfiltr_inst_clk_bfm_clk_clk)        //   clk.clk
	);

initial
begin 
 //fork 
   sin_100();
   sin_50();
   sin_5(); 
 //join_none
#100000000 $stop;
end  
////////////////////////////////////////////////////////////////////
task sin_100(); 
  begin 
  $display ( "begin1" , $time );
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_100;i++)
      begin
        repeat(T_100) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_100_i = mem_100_a[i];    $display ( "begin2" , $time ); end   
  $display ( "begin3" , $time ); 
      end 
  $display ( "begin4" , $time );
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
  $display ( "begin5" , $time );
    for (int i=0;i<K*N_100;i++)
      begin
  $display ( "begin6" , $time );
        repeat(T_100) begin
  $display ( "begin7" , $time );
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
  $display ( "begin8" , $time );
        signal_100_i = mem_100_b[i];   end   
      end 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_100;i++)
      begin
        repeat(T_100) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_100_i = mem_100_c[i];   end   
      end 
  end
endtask 

task sin_50(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_50;i++)
      begin
        repeat(T_50) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_50_i = mem_50_a[i];   end   
      end 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_50;i++)
      begin
        repeat(T_50) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_50_i = mem_50_b[i];   end   
      end 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_50;i++)
      begin
        repeat(T_50) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_50_i = mem_50_c[i];   end   
      end 
  end
endtask 

task sin_5(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_5;i++)
      begin
        repeat(T_5) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_5_i = mem_5_a[i];   end   
      end 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_5;i++)
      begin
        repeat(T_5) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_5_i = mem_5_b[i];   end   
      end 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_5;i++)
      begin
        repeat(T_5) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_5_i = mem_5_c[i];   end   
      end 
  end
endtask 
 
//////////////////////////////////////////////////////////////////////////// /*
/*
task sin_5_a(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_5;i++)
      begin
        repeat(T_5) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_5_i = mem_5_a[i];   end   
      end 
  end
endtask 
///////////////////////////////////////////////////////////////////
task sin_100_b(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_100;i++)
      begin
        repeat(T_100) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_100_i = mem_100_b[i];   end   
      end 
  end
endtask 

task sin_50_b(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_50;i++)
      begin
        repeat(T_50) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_50_i = mem_50_b[i];   end   
      end 
  end
endtask 

task sin_5_b(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_5;i++)
      begin
        repeat(T_5) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_5_i = mem_5_b[i];   end   
      end 
  end
endtask 
/////////////////////////////////////////////////////////////////////
task sin_100_c(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_100;i++)
      begin
        repeat(T_100) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_100_i = mem_100_c[i];   end   
      end 
  end
endtask 

task sin_50_c(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_50;i++)
      begin
        repeat(T_50) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_50_i = mem_50_c[i];   end   
      end 
  end
endtask 

task sin_5_c(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N_5;i++)
      begin
        repeat(T_5) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_5_i = mem_5_c[i];   end   
      end 
  end
endtask 

task fork_100(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk); 
            sin_100_a();
            sin_100_b();
            sin_100_c(); 
  end
endtask 

task fork_50(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);
            sin_50_a();
            sin_50_b();
            sin_50_c(); 
  end
endtask 

task fork_5();
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
            sin_5_a();
            sin_5_b();
            sin_5_c(); 
  end
endtask */
endmodule
