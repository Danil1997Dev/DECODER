// SysFiltr_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module SysFiltr_tb (
	);

	wire    sysfiltr_inst_clk_bfm_clk_clk;       // SysFiltr_inst_clk_bfm:clk -> [SysFiltr_inst:clk_clk, SysFiltr_inst_reset_bfm:clk]
	wire    sysfiltr_inst_reset_bfm_reset_reset; // SysFiltr_inst_reset_bfm:reset -> SysFiltr_inst:reset_reset_n

	SysFiltr sysfiltr_inst (
		.clk_clk                 (sysfiltr_inst_clk_bfm_clk_clk),       //            clk.clk
		.decoder_expend_signal_i (),                                    // decoder_expend.signal_i
		.decoder_expend_indicate (),                                    //               .indicate
		.decoder_expend_work     (),                                    //               .work
		.reset_reset_n           (sysfiltr_inst_reset_bfm_reset_reset)  //          reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sysfiltr_inst_clk_bfm (
		.clk (sysfiltr_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) sysfiltr_inst_reset_bfm (
		.reset (sysfiltr_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (sysfiltr_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
