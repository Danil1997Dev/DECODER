// SysFiltr_IIR_0.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module SysFiltr_IIR_0 (
		input  wire        clk_clk,             //        clk.clk
		input  wire [2:0]  iir_direct_opt_i,    // iir_direct.opt_i
		input  wire [2:0]  iir_direct_opt_o,    //           .opt_o
		input  wire        iir_direct_start,    //           .start
		input  wire        iir_direct_clk_en,   //           .clk_en
		input  wire [31:0] iir_export_i_signal, // iir_export.i_signal
		output wire [31:0] iir_export_o_signal, //           .o_signal
		input  wire        reset_reset_n        //      reset.reset_n
	);

	wire  [31:0] nios_data_master_readdata;                          // mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	wire         nios_data_master_waitrequest;                       // mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	wire         nios_data_master_debugaccess;                       // nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	wire  [13:0] nios_data_master_address;                           // nios:d_address -> mm_interconnect_0:nios_data_master_address
	wire   [3:0] nios_data_master_byteenable;                        // nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	wire         nios_data_master_read;                              // nios:d_read -> mm_interconnect_0:nios_data_master_read
	wire         nios_data_master_write;                             // nios:d_write -> mm_interconnect_0:nios_data_master_write
	wire  [31:0] nios_data_master_writedata;                         // nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	wire  [31:0] nios_instruction_master_readdata;                   // mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	wire         nios_instruction_master_waitrequest;                // mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	wire  [13:0] nios_instruction_master_address;                    // nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	wire         nios_instruction_master_read;                       // nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	wire   [2:0] mm_interconnect_0_iir_avalon_slave_0_address;       // mm_interconnect_0:iir_avalon_slave_0_address -> iir:addres
	wire         mm_interconnect_0_iir_avalon_slave_0_write;         // mm_interconnect_0:iir_avalon_slave_0_write -> iir:enabel
	wire  [31:0] mm_interconnect_0_iir_avalon_slave_0_writedata;     // mm_interconnect_0:iir_avalon_slave_0_writedata -> iir:data
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_readdata;    // nios:debug_mem_slave_readdata -> mm_interconnect_0:nios_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_debug_mem_slave_waitrequest; // nios:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_debug_mem_slave_debugaccess; // mm_interconnect_0:nios_debug_mem_slave_debugaccess -> nios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_debug_mem_slave_address;     // mm_interconnect_0:nios_debug_mem_slave_address -> nios:debug_mem_slave_address
	wire         mm_interconnect_0_nios_debug_mem_slave_read;        // mm_interconnect_0:nios_debug_mem_slave_read -> nios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_debug_mem_slave_byteenable;  // mm_interconnect_0:nios_debug_mem_slave_byteenable -> nios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_debug_mem_slave_write;       // mm_interconnect_0:nios_debug_mem_slave_write -> nios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_writedata;   // mm_interconnect_0:nios_debug_mem_slave_writedata -> nios:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                  // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire   [9:0] mm_interconnect_0_ram_s1_address;                   // mm_interconnect_0:ram_s1_address -> ram:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                // mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	wire         mm_interconnect_0_ram_s1_write;                     // mm_interconnect_0:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                 // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire         mm_interconnect_0_ram_s1_clken;                     // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire  [31:0] nios_irq_irq;                                       // irq_mapper:sender_irq -> nios:irq
	wire         rst_controller_reset_out_reset;                     // rst_controller:reset_out -> [iir:reset_l, irq_mapper:reset, mm_interconnect_0:nios_reset_reset_bridge_in_reset_reset, nios:reset_n, ram:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                 // rst_controller:reset_req -> [nios:reset_req, ram:reset_req, rst_translator:reset_req_in]

	Top #(
		.CLK_REF    (50000000),
		.SAMPL_T    (5000000),
		.FRQ_SIGNAL (800000)
	) iir (
		.clk      (clk_clk),                                        //          clock.clk
		.enabel   (mm_interconnect_0_iir_avalon_slave_0_write),     // avalon_slave_0.write
		.data     (mm_interconnect_0_iir_avalon_slave_0_writedata), //               .writedata
		.addres   (mm_interconnect_0_iir_avalon_slave_0_address),   //               .address
		.reset_l  (~rst_controller_reset_out_reset),                //     reset_sink.reset_n
		.opt_i    (iir_direct_opt_i),                               //         direct.opt_i
		.opt_o    (iir_direct_opt_o),                               //               .opt_o
		.start    (iir_direct_start),                               //               .start
		.clk_en   (iir_direct_clk_en),                              //               .clk_en
		.i_signal (iir_export_i_signal),                            //         export.i_signal
		.o_signal (iir_export_o_signal)                             //               .o_signal
	);

	SysFiltr_IIR_0_nios nios (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_data_master_read),                              //                          .read
		.d_readdata                          (nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_data_master_write),                             //                          .write
		.d_writedata                         (nios_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                   //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	SysFiltr_IIR_0_ram ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	SysFiltr_IIR_0_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                          (clk_clk),                                            //                        clk_0_clk.clk
		.nios_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                     // nios_reset_reset_bridge_in_reset.reset
		.nios_data_master_address               (nios_data_master_address),                           //                 nios_data_master.address
		.nios_data_master_waitrequest           (nios_data_master_waitrequest),                       //                                 .waitrequest
		.nios_data_master_byteenable            (nios_data_master_byteenable),                        //                                 .byteenable
		.nios_data_master_read                  (nios_data_master_read),                              //                                 .read
		.nios_data_master_readdata              (nios_data_master_readdata),                          //                                 .readdata
		.nios_data_master_write                 (nios_data_master_write),                             //                                 .write
		.nios_data_master_writedata             (nios_data_master_writedata),                         //                                 .writedata
		.nios_data_master_debugaccess           (nios_data_master_debugaccess),                       //                                 .debugaccess
		.nios_instruction_master_address        (nios_instruction_master_address),                    //          nios_instruction_master.address
		.nios_instruction_master_waitrequest    (nios_instruction_master_waitrequest),                //                                 .waitrequest
		.nios_instruction_master_read           (nios_instruction_master_read),                       //                                 .read
		.nios_instruction_master_readdata       (nios_instruction_master_readdata),                   //                                 .readdata
		.iir_avalon_slave_0_address             (mm_interconnect_0_iir_avalon_slave_0_address),       //               iir_avalon_slave_0.address
		.iir_avalon_slave_0_write               (mm_interconnect_0_iir_avalon_slave_0_write),         //                                 .write
		.iir_avalon_slave_0_writedata           (mm_interconnect_0_iir_avalon_slave_0_writedata),     //                                 .writedata
		.nios_debug_mem_slave_address           (mm_interconnect_0_nios_debug_mem_slave_address),     //             nios_debug_mem_slave.address
		.nios_debug_mem_slave_write             (mm_interconnect_0_nios_debug_mem_slave_write),       //                                 .write
		.nios_debug_mem_slave_read              (mm_interconnect_0_nios_debug_mem_slave_read),        //                                 .read
		.nios_debug_mem_slave_readdata          (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                                 .readdata
		.nios_debug_mem_slave_writedata         (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                                 .writedata
		.nios_debug_mem_slave_byteenable        (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                                 .byteenable
		.nios_debug_mem_slave_waitrequest       (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                                 .waitrequest
		.nios_debug_mem_slave_debugaccess       (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                                 .debugaccess
		.ram_s1_address                         (mm_interconnect_0_ram_s1_address),                   //                           ram_s1.address
		.ram_s1_write                           (mm_interconnect_0_ram_s1_write),                     //                                 .write
		.ram_s1_readdata                        (mm_interconnect_0_ram_s1_readdata),                  //                                 .readdata
		.ram_s1_writedata                       (mm_interconnect_0_ram_s1_writedata),                 //                                 .writedata
		.ram_s1_byteenable                      (mm_interconnect_0_ram_s1_byteenable),                //                                 .byteenable
		.ram_s1_chipselect                      (mm_interconnect_0_ram_s1_chipselect),                //                                 .chipselect
		.ram_s1_clken                           (mm_interconnect_0_ram_s1_clken)                      //                                 .clken
	);

	SysFiltr_IIR_0_irq_mapper irq_mapper (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (nios_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
