// SysFiltr_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
 

module SysFiltr_tb #(parameter
CLK_PRD = 20,// период тактового сигнала в ns
CLK_REF = 50_000_000,// тактоая частота
CLK_SAMPL = 50_000_000,// честота дискретезации
FRQ = 440_000,// честота сигнала
T=CLK_REF/CLK_SAMPL, // период дискретизации  в тактах
N=CLK_SAMPL/FRQ,// период входного сигнала в тактах
K=350// калчество периодов входного сигнала
)(); 
	logic [31:0] signal_i;
	logic indicate; 
	logic work = 1;

	logic [31:0] mema [0:K*N-1];  
	logic [31:0] memb [0:K*N-1];
	logic [31:0] memc [0:K*N-1]; 

	logic sysfiltr_inst_clk_bfm_clk_clk;       // SysFiltr_inst_clk_bfm:clk -> [SysFiltr_inst:clk_clk, SysFiltr_inst_reset_bfm:clk]
	logic sysfiltr_inst_reset_bfm_reset_reset; // SysFiltr_inst_reset_bfm:reset -> SysFiltr_inst:reset_reset_n

	SysFiltr dut (
		.clk_clk                 (sysfiltr_inst_clk_bfm_clk_clk),       //            clk.clk 
		.decoder_expend_signal_i (signal_i),                                    //               .signal_i
		.decoder_expend_work (work),                                    //               .work
		.decoder_expend_indicate (indicate),                                    //               .indicate
		.reset_reset_n           (sysfiltr_inst_reset_bfm_reset_reset)  //          reset.reset_n
	);
  
	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sysfiltr_inst_clk_bfm (
		.clk (sysfiltr_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) sysfiltr_inst_reset_bfm (
		.reset (sysfiltr_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (sysfiltr_inst_clk_bfm_clk_clk)        //   clk.clk
	);

initial
begin 
 wait (sysfiltr_inst_reset_bfm_reset_reset);
#100000
  sina();
//  #10000 
  sinb(); 
//  #10000
  sinc(); 
  #10000 $stop;
end  

task sina(); 
  begin   
  signal_i = 0; 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);
  signal_i = 0;     
    for (int i=0;i<K*N;i++)
      begin
        repeat(T) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_i = mema[i];   end   
      end 
  end
endtask

task sinb(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N;i++)
      begin
        repeat(T) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_i = memb[i];   end   
      end 
  end
endtask

task sinc(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N;i++)
      begin
        repeat(T) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_i = memc[i];   end   
      end 
  end
endtask 

endmodule
 