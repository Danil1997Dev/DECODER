// SysFiltr_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
 

module SysFiltr_tb #(parameter
CLK_PRD = 20,
T=50_000_000/5_000_000, 
N=5_000_000/440_000,
K=50)();
	logic clk_en,start; 
	logic [31:0] signal_i;
	logic [31:0] i,q; 
	logic valid;

	logic [31:0] mema [0:K*N-1];  
	logic [31:0] memb [0:K*N-1];
	logic [31:0] memc [0:K*N-1]; 

	logic sysfiltr_inst_clk_bfm_clk_clk;       // SysFiltr_inst_clk_bfm:clk -> [SysFiltr_inst:clk_clk, SysFiltr_inst_reset_bfm:clk]
	logic sysfiltr_inst_reset_bfm_reset_reset; // SysFiltr_inst_reset_bfm:reset -> SysFiltr_inst:reset_reset_n

	SysFiltr sysfiltr_inst (
		.clk_clk                       (sysfiltr_inst_clk_bfm_clk_clk),       //                     clk.clk
		.cpu_debug_reset_request_reset (sysfiltr_inst_reset_bfm_reset_reset),                                    // cpu_debug_reset_request.reset
		.decoder_expend_valid          (valid),                                    //          decoder_extend.valid
		.decoder_expend_clk_en         (clk_en),                                    //                        .clk_en
		.decoder_expend_i              (i),                                    //                        .i
		.decoder_expend_q              (q),                                    //                        .q
		.decoder_expend_start          (start),                                    //                        .start
		.decoder_expend_signal_i       (signal_i),                                    //                        .signal_i
		.reset_reset_n                 (sysfiltr_inst_reset_bfm_reset_reset)  //                   reset.reset_n
	);
  
	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sysfiltr_inst_clk_bfm (
		.clk (sysfiltr_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) sysfiltr_inst_reset_bfm (
		.reset (sysfiltr_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (sysfiltr_inst_clk_bfm_clk_clk)        //   clk.clk
	);

initial
begin
  #100000
  sina();
//  #10000 
  sinb(); 
//  #10000
  sinc(); 
  #10000 $stop;
end  

task sina(); 
  begin  
  start = 0;
  clk_en = 0;
  signal_i = 0; 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);
  signal_i = 0;   
  start = 1;
  clk_en = 1; 
    for (int i=0;i<K*N;i++)
      begin
        repeat(T) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk); 
        enabel = 1;
        signal_i = mema[i];   end   
      end 
  end
endtask

task sinb(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N;i++)
      begin
        repeat(T) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_i = memb[i];   end   
      end 
  end
endtask

task sinc(); 
  begin 
  @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
    for (int i=0;i<K*N;i++)
      begin
        repeat(T) begin
        @(posedge sysfiltr_inst_clk_bfm_clk_clk);  
        signal_i = memc[i];   end   
      end 
  end
endtask 

endmodule
 